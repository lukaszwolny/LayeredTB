///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//Layerd TB
//EDA
//https://www.edaplayground.com/x/Dsjy
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
`include "interface.sv"
`include "test.sv"
module testbench_top;
  bit clk;
//   bit rst;
  
  //clock generation
  always #5 clk = ~clk;
  
  //interface
  acc_if intf(clk);//, rst
  
  initial
  begin
 	clk = 0;
  end
  
  //testcase
  test test1(intf);
  
  //DUT
  accumulator #(
    .WIDTH(8)
  ) u_acc (
    .clk(intf.clk),
    .rst(intf.rst),
    .in(intf.in),
    .ceAcu(intf.ceAcu),
    .out(intf.out)
  );
  
  initial
  begin 
    $dumpfile("dump.vcd"); $dumpvars;
  end
endmodule
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////